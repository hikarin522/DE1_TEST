
module CLOCK24(
	input CLOCK_50,
	input [3:0] KEY,
	output [9:0] LEDR,
	output [6:0] HEX0, HEX1, HEX2, HEX3, HEX4, HEX5
);

_CLOCK24 _CLOCK24(CLOCK_50, 1'b0, KEY[2:0], LEDR, HEX0, HEX1, HEX2, HEX3, HEX4, HEX5);

endmodule

module _CLOCK24(
	input CLK, RST,
	input [2:0] nBUTTON,
	output [9:0] LEDR,
	output [6:0] nHEX0, nHEX1, nHEX2, nHEX3, nHEX4, nHEX5
);

wire CASEC, CAMIN;
wire MODE, SELECT, ADJUST;
wire SECCLR, MININC, HOURINC;
wire SECON, MINON, HOURON;
wire EN1HZ, SIG2HZ;
wire [2:0] btn;
wire [3:0] SECL, MINL, HOURL;
wire [2:0] SECH, MINH;
wire [1:0] HOURH;

CNT1SEC CNT1SEC(CLK, RST, EN1HZ, SIG2HZ);
BTN_IN BTN_IN(.CLK(CLK), .RST(RST), .nBIN(nBUTTON), .BOUT({MODE, SELECT, ADJUST}));
SECCNT SEC(CLK, RST, EN1HZ, SECCLR, SECH, SECL, CASEC);
MINCNT MIN(CLK, RST, CASEC, MININC, MINH, MINL, CAMIN);
HOURCNT HOUR(CLK, RST, CAMIN, HOURINC, HOURH, HOURL);
STATE STATE(CLK, RST, SIG2HZ, MODE, SELECT, ADJUST, SECCLR, MININC, HOURINC, SECON, MINON, HOURON);
SEG7DEC SL(SECL, SECON, nHEX0);
SEG7DEC SH({1'b0, SECH}, SECON, nHEX1);
SEG7DEC ML(MINL, MINON, nHEX2);
SEG7DEC MH({1'b0, MINH}, MINON, nHEX3);
SEG7DEC HL(HOURL, HOURON, nHEX4);
SEG7DEC HH({2'b00, HOURH}, HOURON, nHEX5);

assign LEDR[3:0] = (SECON == 1'b1) ? SECL : 4'h0;
assign LEDR[6:4] = (SECON == 1'b1) ? SECH : 3'h0;
assign LEDR[9:7] = 3'h0;

endmodule
